library ieee;
use ieee.std_logic_1164.all;

package mux_p is
  type slv_array_t is array (natural range <>) of std_logic_vector (4 downto 0);
end package;

package body mux_p is
end package body;